
---------------------------------------------------------------------------------
-- Univ. of Chicago  
--    
--
-- PROJECT:      ANNIE - ACDC
-- FILE:         trigger.vhd
-- AUTHOR:       D. Greenshields
-- DATE:         May 2021
--
-- DESCRIPTION:  trigger processes
---------------------------------------------------------------------------------

	
library IEEE;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;
use work.defs.all;
use work.LibDG.pulseSync;
use work.LibDG.pulseSync2;
use work.LibDG.manchester_decoder;
use work.components.all;

entity trigger is
	port(
			clock			 : in	clock_type;
			reset			 : in	reset_type;   
			systemTime		 : in  std_logic_vector(63 downto 0);
            wrTime_pps       : in std_logic_vector(31 downto 0);
            wrTime_fast      : in std_logic_vector(31 downto 0);
			trigSetup		 : in	trig_type;
			selfTrig		 : in 	selfTrig_type;
			trigInfo		 : out	trigInfo_type;
			acc_trig		 : in	std_logic;	-- trig from central card (LVDS)
			self_trig		 : in	std_logic;	
			digitize_request : out	std_logic;
			digitize_done	 : in	std_logic;
			eventCount		 : out	std_logic_vector(31 downto 0);
			sys_timestamp	 : out std_logic_vector(63 downto 0);
            sys_ts_read      : in std_logic;
            sys_ts_valid     : out std_logic;
            wr_timestamp	 : out std_logic_vector(63 downto 0);
            wr_ts_read       : in std_logic;
            wr_ts_valid      : out std_logic;
            backpressure_in  : in std_logic;
            backpressure_in_acdc : in std_logic;
			busy			 : out std_logic;
			trig_clear		 : buffer std_logic;
			trig_out		 : buffer std_logic;
            trig_out_debug   : out std_logic;
			trig_count_all   : out std_logic_vector(15 downto 0);
            trig_count	     : out std_logic_vector(15 downto 0);
            trig_count_reset : in  std_logic;
            wr_timeOcc       : out std_logic_vector(3 downto 0);
            sys_timeOcc      : out std_logic_vector(3 downto 0)
			);
end trigger;

architecture vhdl of trigger is

    signal 	acc_trig_in:	std_logic;
  	signal 	acc_trig_in_x:	std_logic;
	signal 	trig_latch:	std_logic;
	signal 	trig_latch_x:	std_logic;
	signal 	trig_latch_z:	std_logic;
	signal 	trig_latch_z2:	std_logic;
    signal 	trig_latch_z3:	std_logic;
    signal  wr_trig_z1 : std_logic;
    signal  wr_trig_z2 : std_logic;
    signal  wr_trig_z3 : std_logic;
	signal	trig_common: std_logic;
	signal	timestamp_z: std_logic_vector(63 downto 0);
    signal	timestamp_z2: std_logic_vector(63 downto 0);
    signal  wrTime_pps_z   : std_logic_vector(31 downto 0);
    signal  wrTime_fast_z  : std_logic_vector(31 downto 0);
	signal	prev_mode: natural;
	signal 	acc_trig_x:	std_logic;
	signal	mode_z: natural;
    signal  save_timestamps : std_logic;
    signal  save_timestamps_wr_sync : std_logic;
    signal  save_timestamps_sys_sync : std_logic;
    signal  wr_ts_fifo_empty : std_logic;
    signal  sys_ts_fifo_empty : std_logic;
	
begin  



-- brief description:
---------------------
-- A trigger is detected which has different sources depending on the mode:-
--
-- sma input
-- acc (sma, software or pps)
-- self trigger (generated by psec4 chips when signal level exceeds threshold on selected channels
--
-- For some modes a validation signal must also be received within a certain time of the trigger
-- This can come from sma input or acc
--



---------------------------------------
-- TRIGGER SELECT
---------------------------------------

-- decode acc_trig
manchester_decoder_inst: manchester_decoder
  port map (
    clk    => clock.x8,
    resetn => not reset.global,
    i      => acc_trig,
    q      => acc_trig_in);

trig_out_debug <= acc_trig_in;

TRIG_ACCEPT_SEL: process(all)
begin
    case trigSetup.mode is
        when 0 => trig_common <= '0';          -- mode 0 trigger off
        when 1 => trig_common <= acc_trig_in;  -- mode 1 external source
        when 2 => trig_common <= self_trig;    -- mode 2 self trigger
        when 3 => trig_common <= self_trig;    -- mode 3 self trigger with ACC accept
        when others => trig_common <= '0';
    end case;
end process;

---------------------------------------
-- TRIGGER LATCH
---------------------------------------


-- Edge detect
TRIG_EDGE_DETECT: process(trig_common, trig_clear, reset.global)
begin
	if (trig_clear = '1' or reset.global = '1') then
		trig_latch <= '0';
	elsif (rising_edge(trig_common)) then
		trig_latch <= '1';
	end if;
end process;

trig_out <= trig_latch;			-- trigger to PSEC chips


---------------------------------------
-- TRIGGER TIMESTAMP GENERATOR
---------------------------------------
-- generate a timestamp value for when the trigger latch goes high 

TIMESTAMP_GEN: process(clock.x8)
begin
	if (rising_edge(clock.x8)) then
		trig_latch_z <= trig_latch;		-- synchronize to fast clock
		trig_latch_z2 <= trig_latch_z;
        trig_latch_z3 <= trig_latch_z2;
		if (trig_latch_z2 = '1' and trig_latch_z3 = '0') then	-- rising edge
			timestamp_z <= systemTime;
		end if;
	end if;
end process;

pulseSync2_sys_timesave: pulseSync2
  port map (
    src_clk      => clock.sys,
    src_pulse    => save_timestamps,
    src_aresetn  => not reset.global,
    dest_clk     => clock.x4,
    dest_pulse   => save_timestamps_sys_sync,
    dest_aresetn => not reset.global);

sys_ts_valid <= not sys_ts_fifo_empty;

-- Cyclone IV FIFO cannot be clocked at 320 MHz, so lets bring the data to the
-- 160 MHz domain first (should have plenty of time, from state machine delay
-- and trigger sync stages above)
time_SYS_slowdown : process(clock.x4)
begin
  if rising_edge(clock.x4) then
    timestamp_z2 <= timestamp_z;
  end if;
end process;

timeFifo_SYS: timeFifo
  port map (
    aclr    => reset.global,
    wrclk   => clock.x4,
    wrreq   => save_timestamps_sys_sync,
    data    => timestamp_z2,
    wrfull  => open,
    
    rdclk   => clock.serial25,
    rdreq   => sys_ts_read,
    q       => sys_timestamp,
    rdempty => sys_ts_fifo_empty,
    rdusedw => sys_timeOcc
    );

WR_TIMESTAMP_GEN: process(clock.wr250)
begin
  if (rising_edge(clock.wr250)) then
    wr_trig_z1 <= trig_latch;		-- synchronize to fast clock
    wr_trig_z2 <= wr_trig_z1;
    wr_trig_z3 <= wr_trig_z2;
    if (wr_trig_z2 = '1' and wr_trig_z3 = '0') then	-- rising edge
      wrTime_pps_z  <= wrTime_pps; 
      wrTime_fast_z <= wrTime_fast; 
    end if;
  end if;
end process;

pulseSync2_wr_timesave: pulseSync2
  port map (
    src_clk      => clock.sys,
    src_pulse    => save_timestamps,
    src_aresetn  => not reset.global,
    dest_clk     => clock.wr250,
    dest_pulse   => save_timestamps_wr_sync,
    dest_aresetn => not reset.wr);

-- hack to keep fifo "open" if clock is not present
wr_ts_valid <= (not wr_ts_fifo_empty) or (not clock.wrpllLock);

timeFifo_WR: timeFifo
  port map (
    aclr    => reset.wr,
    wrclk   => clock.wr250,
    wrreq   => save_timestamps_wr_sync,
    data    => wrTime_pps_z & wrTime_fast_z,
    wrfull  => open,
    
    rdclk   => clock.serial25,
    rdreq   => wr_ts_read,
    q       => wr_timestamp,
    rdempty => wr_ts_fifo_empty,
    rdusedw => wr_timeOcc
    );

	
---------------------------------------
-- TRIGGER CONTROL STATE MACHINE
---------------------------------------

TRIG_CTRL: process(clock.sys)

type state_type is (
	TRIG_RESET, 
	TRIG_WAIT, 
	TRIG_CONFIRM,
	DIGITIZE_INIT, 
	DIGITIZE_WAIT, 
	TRIG_DONE
);
	
variable t: natural range 0 to 127;
variable state: state_type;

begin
	if (rising_edge(clock.sys)) then
	
		-- synchronize to sys clock
		trig_latch_x <= trig_latch;
        acc_trig_in_x <= acc_trig_in;
		
		-- reset trigger state if mode change
		prev_mode <= trigSetup.mode;
		if (prev_mode /= trigSetup.mode or trigSetup.resetReq = '1') then 
			state := TRIG_RESET; 
		end if;			
				
		-- global reset or event count reset request
		if (reset.global = '1' or trigSetup.eventAndTime_reset = '1') then 

            digitize_request <= '0';
			state := TRIG_RESET;
			eventCount <= X"00000000";
            save_timestamps <= '0';
            trig_count_all  <= (others => '0');
            trig_count	    <= (others => '0');

		else
		
			case state is
			
				when TRIG_RESET =>
				
					trig_clear <= '1';		-- clear the latches
					if (trig_latch_x = '0') then state := TRIG_WAIT; end if;		-- verify the latch is clear before waiting for a latch high signal
	
	
				when TRIG_WAIT =>				-- wait for an incoming trigger trigger signal
									
                    trig_clear <= '0';		-- enable the trigger latches
                    save_timestamps <= '0';

                    t := trigSetup.timeout;
                    
					if (trig_latch_x = '1') then		-- trigger latch went high					
                      state := TRIG_CONFIRM;
                      trig_count_all <= std_logic_vector(unsigned(trig_count_all) + 1);
					end if;
				
						
				when TRIG_CONFIRM =>				-- timestamp value has already been latched but copy its value and sync to sys clk

                    t := t;
                    save_timestamps <= '0';
                    
                    if backpressure_in = '1' or backpressure_in_acdc = '1' then
                      state := TRIG_RESET;
                    else
                      case trigSetup.mode is
                        when 0 => state := TRIG_RESET;     -- mode 0 trigger off
                        when 1 => state := DIGITIZE_INIT;  -- mode 1 external source
                        when 2 => state := DIGITIZE_INIT;  -- mode 2 self trigger
                        when 3 =>                          -- mode 3 self trigger with ACC accept
                          if acc_trig_in_x = '1' then
                            state := DIGITIZE_INIT;
                          elsif t = 0 then
                            state := TRIG_RESET;
                          else
                            state := state;
                            t := t - 1;
                          end if;
                          
                        when others => state := TRIG_RESET;
                      end case;
                    end if;

                    
				when DIGITIZE_INIT =>				-- request to start transfer of data from psec to fpga

                    save_timestamps <= '1';
                    
                    trig_count <= std_logic_vector(unsigned(trig_count) + 1);
                  
					digitize_request <= '1';
					state := DIGITIZE_WAIT;
				
				
				when DIGITIZE_WAIT =>				-- wait for the PSEC chip data to be transferred to the fpga RAM

                    save_timestamps <= '0';
                  
					digitize_request <= '0';
					if (digitize_done = '1') then state := TRIG_DONE; end if;
				
				
				when TRIG_DONE =>

                    eventCount <= eventCount + 1;
					state := TRIG_RESET;
					
			end case;
				
			if (state = TRIG_WAIT) then busy <= '0'; else busy <= '1'; end if;
		
		end if;
		
	end if;
	
end process;


--
--trigInfo(0,0) <= beamgate_timestamp(63 downto 48);
--trigInfo(0,1) <= beamgate_timestamp(47 downto 32);
--trigInfo(0,2) <= beamgate_timestamp(31 downto 16);
--trigInfo(0,3) <= beamgate_timestamp(15 downto 0);

trigInfo(0,4)(15 downto 12) <= std_logic_vector(to_unsigned(trigSetup.mode, 4));
trigInfo(0,4)(11 downto 10) <= trigSetup.sma_invert & selfTrig.sign;
trigInfo(0,4)(9 downto 0) <= "00000" & std_logic_vector(to_unsigned(selfTrig.coincidence_min, 5));

--
trigInfo(1,0) <= "0000000000" & selfTrig.mask(0);
trigInfo(1,1) <= "0000000000" & selfTrig.mask(1);
trigInfo(1,2) <= "0000000000" & selfTrig.mask(2);
trigInfo(1,3) <= "0000000000" & selfTrig.mask(3);
trigInfo(1,4) <= "0000000000" & selfTrig.mask(4);

--
trigInfo(2,0) <= x"0" & std_logic_vector(to_unsigned(selfTrig.threshold(0, 0), 12));
trigInfo(2,1) <= x"0" & std_logic_vector(to_unsigned(selfTrig.threshold(1, 0), 12));
trigInfo(2,2) <= x"0" & std_logic_vector(to_unsigned(selfTrig.threshold(2, 0), 12));
trigInfo(2,3) <= x"0" & std_logic_vector(to_unsigned(selfTrig.threshold(3, 0), 12));
trigInfo(2,4) <= x"0" & std_logic_vector(to_unsigned(selfTrig.threshold(4, 0), 12));



------------------------------
-- TRIGGER RATE COUNTER
------------------------------
-- count the number of trig events in one second 

--RATE_COUNT_GEN: process(clock.sys)
--variable count: natural;
--variable t: natural;
--begin
--	if (rising_edge(clock.sys)) then
--		
--		if (reset.global = '1' or trigSetup.eventAndTime_reset = '1') then
--		
--			t := 0;
--			count := 0;
--			trig_rate_count <= 0;
--			
--			
--		else
--		
--		
--			if (trig_event = '1') then
--				if (count < trigRate_MaxCount) then count := count + 1; end if;
--			end if;				
--			
--			t := t + 1;		-- clock cycle counter
--			 
--			if (t = 40000000) then		-- after 1 second record the count and then reset 
--
--				t := 0;
--				trig_rate_count <= count;
--				count := 0;
--				
--			end if;
--			
--		end if;
--		
--	end if;
--end process;

	
end vhdl;






